module tile_map ( output logic [0:29][0:39] tile );
	always_comb
	begin
		tile =
		{
			40'h0, // will occupy about two line if not zero. HOW COME?!!!!
			40'h8000000001, // 1
			40'h8000000001, // 2
			40'h8000000001, // 3
			40'h81FF000001, // 4
			40'h8003000001, // 5
			40'h8000FFFFFF, // 6
			40'h8000000001, // 7
			40'hFF00000001, // 8
			40'h8000000001, // 9
			40'h8000000001, // 10
			40'h8000000001, // 11
			40'hFFFFFFFFE1, // 12
			40'h80000003E1, // 13
			40'h8000000001, // 14
			40'h800000000F, // 15
			40'h80FFFFF001, // 16
			40'h8000003FFF, // 17
			40'h8000000001, // 18
			40'hF000000001, // 19
			40'h8000000001, // 20
			40'hFFFFF80001, // 21
			40'h8000008001, // 22
			40'h800000FFC1, // 23
			40'h8000000001, // 24
			40'hFFFF000001, // 25
			40'h800000000F, // 26
			40'h8000000001, // 27
			40'h8000000001, // 28
			40'hFFFFFFFFFF  // 29
		};
	end
					
endmodule
